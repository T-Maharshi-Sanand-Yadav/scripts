`timescale 1ns / 1ps
module nor_gate_level_modelling(y,a,b);
output y;
input a,b;
nor x1(y,a,b);
endmodule
