************************************************************************
* auCdl Netlist:
* 
* Library Name:  exnor_gate
* Top Cell Name: exnor
* View Name:     schematic
* Netlisted on:  Mar  1 23:01:22 2023
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: inverter
* Cell Name:    inverter
* View Name:    schematic
************************************************************************
simulator lang=spice
.SUBCKT inverter A GND VDD Y
*.PININFO A:I Y:O GND:B VDD:B
MNM0 Y A GND GND nmos W=2u L=180n M=1
MPM0 Y A VDD VDD pmos W=2u L=180n M=1
.ENDS

************************************************************************
* Library Name: exor_gate
* Cell Name:    exor
* View Name:    schematic
************************************************************************

.SUBCKT exor a b gnd vdd Y
*.PININFO a:I b:I Y:O gnd:B vdd:B
MPM5 Y b net23 vdd pmos W=2u L=180n M=1
MPM4 net23 abar vdd vdd pmos W=2u L=180n M=1
MPM1 Y bbar net24 vdd pmos W=2u L=180n M=1
MPM0 net24 a vdd vdd pmos W=2u L=180n M=1
MNM3 net21 bbar gnd gnd nmos W=2u L=180n M=1
MNM2 Y abar net21 gnd nmos W=2u L=180n M=1
MNM1 net22 b gnd gnd nmos W=2u L=180n M=1
MNM0 Y a net22 gnd nmos W=2u L=180n M=1
XI1 a gnd vdd abar / inverter
XI0 b gnd vdd bbar / inverter
.ENDS

************************************************************************
* Library Name: exnor_gate
* Cell Name:    exnor
* View Name:    schematic
************************************************************************

.SUBCKT exnor A B GND VDD Y
*.PININFO A:I B:I Y:O GND:B VDD:B
XI0 A B GND VDD net14 / exor
XI1 net14 GND VDD Y / inverter
.ENDS

