************************************************************************
* auCdl Netlist:
* 
* Library Name:  inverter
* Top Cell Name: inverter
* View Name:     schematic
* Netlisted on:  Mar  2 02:32:26 2023
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: inverter
* Cell Name:    inverter
* View Name:    schematic
************************************************************************

.SUBCKT inverter A GND VDD Y
*.PININFO A:I Y:O GND:B VDD:B
MNM0 Y A GND GND g45n1svt m=1 l=45n w=120n
MPM0 Y A VDD VDD g45p1svt m=1 l=45n w=120n
.ENDS

