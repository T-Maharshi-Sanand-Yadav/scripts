`timescale 1ns / 1ps
module not_gate_level_modelling(y,a);
output y;
input a;
not x1(y,a);
endmodule

