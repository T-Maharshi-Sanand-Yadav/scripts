************************************************************************
* auCdl Netlist:
* 
* Library Name:  or_gate
* Top Cell Name: or
* View Name:     schematic
* Netlisted on:  Mar  1 23:49:45 2023
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: nor_gate
* Cell Name:    nor
* View Name:    schematic
************************************************************************
simulator lang=spice
.SUBCKT nor A B GND VDD Y
*.PININFO A:I B:I Y:O GND:B VDD:B
MNM1 Y B GND GND nmos W=2u L=180n M=1
MNM0 Y A GND GND nmos W=2u L=180n M=1
MPM1 net18 A VDD VDD pmos W=2u L=180n M=1
MPM0 Y B net18 VDD pmos W=2u L=180n M=1
.ENDS

************************************************************************
* Library Name: inverter
* Cell Name:    inverter
* View Name:    schematic
************************************************************************

.SUBCKT inverter A GND VDD Y
*.PININFO A:I Y:O GND:B VDD:B
MNM0 Y A GND GND nmos W=2u L=180n M=1
MPM0 Y A VDD VDD pmos W=2u L=180n M=1
.ENDS

************************************************************************
* Library Name: or_gate
* Cell Name:    or
* View Name:    schematic
************************************************************************

.SUBCKT or A B GND VDD Y
*.PININFO A:I B:I Y:O GND:B VDD:B
XI0 A B GND VDD net14 / nor
XI1 net14 GND VDD Y / inverter
.ENDS

