`timescale 1ns / 1ps
module or_gate_level_modelling(y,a,b);
output y;
input a,b;
or x1(y,a,b);
endmodule

