************************************************************************
* auCdl Netlist:
* 
* Library Name:  nand_gate
* Top Cell Name: nand
* View Name:     schematic
* Netlisted on:  Mar  1 23:47:43 2023
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: nand_gate
* Cell Name:    nand
* View Name:    schematic
************************************************************************
simulator lang=spice
.SUBCKT nand A B GND VDD Y
*.PININFO A:I B:I Y:O GND:B VDD:B
MNM1 net20 B GND GND nmos W=2u L=180n M=1
MNM0 Y A net20 GND nmos W=2u L=180n M=1
MPM1 Y B VDD VDD pmos W=2u L=180n M=1
MPM0 Y A VDD VDD pmos W=2u L=180n M=1
.ENDS

