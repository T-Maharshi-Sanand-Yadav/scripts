************************************************************************
* auCdl Netlist:
* 
* Library Name:  invert
* Top Cell Name: inv
* View Name:     schematic
* Netlisted on:  Mar  1 23:55:38 2023
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: invert
* Cell Name:    inv
* View Name:    schematic
************************************************************************

.SUBCKT inv a gnd vdd y
*.PININFO a:I y:O gnd:B vdd:B
MNM0 y a gnd gnd nmos1v m=1 l=100n w=120n
MPM0 y a vdd vdd pmos1v m=1 l=100n w=360n
.ENDS

