`timescale 1ns / 1ps
module not_data_flow_modelling(y,a);
output y;
input a;
assign y = ~a;
endmodule

