`timescale 1ns / 1ps
module xor_gate_level_modelling(y,a,b);
output y;
input a,b;
xor x1(y,a,b);
endmodule
