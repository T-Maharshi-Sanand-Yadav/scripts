************************************************************************
* auCdl Netlist:
* 
* Library Name:  or_gate
* Top Cell Name: or
* View Name:     schematic
* Netlisted on:  Mar  1 23:57:37 2023
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: nor_gate
* Cell Name:    nor
* View Name:    schematic
************************************************************************

.SUBCKT nor a b gnd vdd y
*.PININFO a:I b:I y:O gnd:B vdd:B
MNM1 y b gnd gnd nmos1v m=1 l=100n w=120n
MNM0 y a gnd gnd nmos1v m=1 l=100n w=120n
MPM1 y b net18 vdd pmos1v m=1 l=100n w=360n
MPM0 net18 a vdd vdd pmos1v m=1 l=100n w=360n
.ENDS

************************************************************************
* Library Name: invert
* Cell Name:    inv
* View Name:    schematic
************************************************************************

.SUBCKT inv a gnd vdd y
*.PININFO a:I y:O gnd:B vdd:B
MNM0 y a gnd gnd nmos1v m=1 l=100n w=120n
MPM0 y a vdd vdd pmos1v m=1 l=100n w=360n
.ENDS

************************************************************************
* Library Name: or_gate
* Cell Name:    or
* View Name:    schematic
************************************************************************

.SUBCKT or a b gnd vdd y
*.PININFO a:I b:I y:O gnd:B vdd:B
XI0 a b gnd vdd net13 / nor
XI1 net13 gnd vdd y / inv
.ENDS

