************************************************************************
* auCdl Netlist:
* 
* Library Name:  nor_gate
* Top Cell Name: nor
* View Name:     schematic
* Netlisted on:  Mar  1 23:48:13 2023
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: nor_gate
* Cell Name:    nor
* View Name:    schematic
************************************************************************
simulator lang=spice
.SUBCKT nor A B GND VDD Y
*.PININFO A:I B:I Y:O GND:B VDD:B
MNM1 Y B GND GND nmos W=2u L=180n M=1
MNM0 Y A GND GND nmos W=2u L=180n M=1
MPM1 net18 A VDD VDD pmos W=2u L=180n M=1
MPM0 Y B net18 VDD pmos W=2u L=180n M=1
.ENDS

