************************************************************************
* auCdl Netlist:
* 
* Library Name:  nor_gate
* Top Cell Name: nor
* View Name:     schematic
* Netlisted on:  Mar  1 23:56:45 2023
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: nor_gate
* Cell Name:    nor
* View Name:    schematic
************************************************************************

.SUBCKT nor a b gnd vdd y
*.PININFO a:I b:I y:O gnd:B vdd:B
MNM1 y b gnd gnd nmos1v m=1 l=100n w=120n
MNM0 y a gnd gnd nmos1v m=1 l=100n w=120n
MPM1 y b net18 vdd pmos1v m=1 l=100n w=360n
MPM0 net18 a vdd vdd pmos1v m=1 l=100n w=360n
.ENDS

