************************************************************************
* auCdl Netlist:
* 
* Library Name:  and_gate
* Top Cell Name: and
* View Name:     schematic
* Netlisted on:  Mar  1 23:00:46 2023
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: nand_gate
* Cell Name:    nand
* View Name:    schematic
************************************************************************
simulator lang=spice
.SUBCKT nand A B GND VDD Y
*.PININFO A:I B:I Y:O GND:B VDD:B
MNM1 net20 B GND GND nmos W=2u L=180n M=1
MNM0 Y A net20 GND nmos W=2u L=180n M=1
MPM1 Y B VDD VDD pmos W=2u L=180n M=1
MPM0 Y A VDD VDD pmos W=2u L=180n M=1
.ENDS

************************************************************************
* Library Name: inverter
* Cell Name:    inverter
* View Name:    schematic
************************************************************************

.SUBCKT inverter A GND VDD Y
*.PININFO A:I Y:O GND:B VDD:B
MNM0 Y A GND GND nmos W=2u L=180n M=1
MPM0 Y A VDD VDD pmos W=2u L=180n M=1
.ENDS

************************************************************************
* Library Name: and_gate
* Cell Name:    and
* View Name:    schematic
************************************************************************

.SUBCKT and A B GND VDD Y
*.PININFO A:I B:I Y:O GND:B VDD:B
XI0 A B GND VDD net15 / nand
XI1 net15 GND VDD Y / inverter
.ENDS

