************************************************************************
* auCdl Netlist:
* 
* Library Name:  nor_gate
* Top Cell Name: nor
* View Name:     schematic
* Netlisted on:  Mar  2 02:33:21 2023
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: nor_gate
* Cell Name:    nor
* View Name:    schematic
************************************************************************

.SUBCKT nor A B GND VDD Y
*.PININFO A:I B:I Y:O GND:B VDD:B
MNM1 Y B GND GND g45n1svt m=1 l=45n w=120n
MNM0 Y A GND GND g45n1svt m=1 l=45n w=120n
MPM1 net17 A VDD VDD g45p1svt m=1 l=45n w=120n
MPM0 Y B net17 VDD g45p1svt m=1 l=45n w=120n
.ENDS

