`timescale 1ns / 1ps
module and_gate_level_modelling(y,a,b);
output y;
input a,b;
and x1(y,a,b);
endmodule


